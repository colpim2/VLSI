library ieee;
use ieee.std_logic_1164.all;

entity conta3display is
port(clk: in std_logic;
	  ssg0: out std_logic_vector(6 downto 0);
	  ssg1: out std_logic_vector(6 downto 0);
	  ssg2: out std_logic_vector(6 downto 0));
end entity;

architecture a of conta3display is

signal bandera, bandera2: std_logic;
signal banderaSal, banderaSal2: std_logic;
signal conteo, conteo2: integer range 0 to 9;

begin
	
	u4: entity work.contador(arqcontador)  port map(clk, ssg0, bandera);
	u5: entity work.cont(arqcont) 			port map(bandera, conteo, banderaSal);
	u6: entity work.ss7(arqss7)   			port map(conteo, ssg1);
	u7: entity work.cont(arqcont) 			port map(banderaSal, conteo2, banderaSal2);
	u8: entity work.ss7(arqss7)   			port map(conteo2, ssg2);
	
end architecture;