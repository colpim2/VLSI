library ieee;
use ieee.std_logic_1164.all;

entity cont is
port(clk: in std_logic;
	  reset: in std_logic);
end entity;

architecture arqcontr of cont is

signal clkl: std_logic;
signal a: integer range 0 to 9;

begin
	
end architecture;